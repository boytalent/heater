module lfsr_checker(
    input   logic           clk,
    input   logic           reset,
    input   logic   [31:0]  datain,
    output  logic           error);

    logic   [31:0]  next_lfsr, next_lfsr_q;

    lfsr #(.WIDTH(32)) lfsr_inst (.datain(datain), .dataout(next_lfsr));

    always_ff @(posedge clk) next_lfsr_q <= next_lfsr;
    logic compare;
    always_ff @(posedge clk) if (next_lfsr_q == datain) compare <= 1; else compare <= 0;
    always_ff @(posedge clk) if (reset == 1) error <= 0; else if (!compare) error <= 1;

endmodule

